module greensc (
  input [7:0] in_r,
  input [7:0] in_g,
  input [7:0] in_b,
  
  output [7:0] out_r,
  output [7:0] out_g,
  output [7:0] out_b
);
  
  
endmodule
