module gauss(
input clk,
input [7:0] r, b , g,
input [12:0] col,
input wr_en,
input filt_sel,
output [7:0] out_r, out_g, out_b

);
//
//saturate satr(.in(r10_out[0][17:8]), .out(out_r));
//saturate satb(.in(tmp_1[1][17:8]), .out(out_g));
//saturate satg(.in(tmp_1[2][17:8]), .out(out_b));
wire [7:0] gauss_r, gauss_g, gauss_b;
wire [7:0] r0_out, r1_out, r2_out, r3_out, r4_out, r5_out, r6_out, r7_out, r8_out, r9_out, r10_out;
wire [7:0] g0_out, g1_out, g2_out, g3_out, g4_out, g5_out, g6_out, g7_out, g8_out, g9_out, g10_out;
wire [7:0] b0_out, b1_out, b2_out, b3_out, b4_out, b5_out, b6_out, b7_out, b8_out, b9_out, b10_out;

assign out_r = r10_out;
assign out_g = g10_out;
assign out_b = b10_out;
ram r0(.clk(clk), .wr_en(wr_en), .addr(col), .data_in(r), .data_out(r0_out));
ram r1(.clk(clk), .wr_en(wr_en), .addr(col + 1), .data_in(r0_out), .data_out(r1_out));
ram r2(.clk(clk), .wr_en(wr_en), .addr(col + 2), .data_in(r1_out), .data_out(r2_out));
ram r3(.clk(clk), .wr_en(wr_en), .addr(col + 3), .data_in(r2_out), .data_out(r3_out));
ram r4(.clk(clk), .wr_en(wr_en), .addr(col + 4), .data_in(r3_out), .data_out(r4_out));
ram r5(.clk(clk), .wr_en(wr_en), .addr(col + 5), .data_in(r4_out), .data_out(r5_out));
ram r6(.clk(clk), .wr_en(wr_en), .addr(col + 6), .data_in(r5_out), .data_out(r6_out));
ram r7(.clk(clk), .wr_en(wr_en), .addr(col + 7), .data_in(r6_out), .data_out(r7_out));
ram r8(.clk(clk), .wr_en(wr_en), .addr(col + 8), .data_in(r7_out), .data_out(r8_out));
ram r9(.clk(clk), .wr_en(wr_en), .addr(col + 9), .data_in(r8_out), .data_out(r9_out));
ram r10(.clk(clk), .wr_en(wr_en), .addr(col + 10), .data_in(r9_out), .data_out(r10_out));

ram g0(.clk(clk), .wr_en(wr_en), .addr(col), .data_in(r), .data_out(g0_out));
ram g1(.clk(clk), .wr_en(wr_en), .addr(col + 1), .data_in(g0_out), .data_out(g1_out));
ram g2(.clk(clk), .wr_en(wr_en), .addr(col + 2), .data_in(g1_out), .data_out(g2_out));
ram g3(.clk(clk), .wr_en(wr_en), .addr(col + 3), .data_in(g2_out), .data_out(g3_out));
ram g4(.clk(clk), .wr_en(wr_en), .addr(col + 4), .data_in(g3_out), .data_out(g4_out));
ram g5(.clk(clk), .wr_en(wr_en), .addr(col + 5), .data_in(g4_out), .data_out(g5_out));
ram g6(.clk(clk), .wr_en(wr_en), .addr(col + 6), .data_in(g5_out), .data_out(g6_out));
ram g7(.clk(clk), .wr_en(wr_en), .addr(col + 7), .data_in(g6_out), .data_out(g7_out));
ram g8(.clk(clk), .wr_en(wr_en), .addr(col + 8), .data_in(g7_out), .data_out(g8_out));
ram g9(.clk(clk), .wr_en(wr_en), .addr(col + 9), .data_in(g8_out), .data_out(g9_out));
ram g10(.clk(clk), .wr_en(wr_en), .addr(col + 10), .data_in(r9_out), .data_out(g10_out));

ram b0(.clk(clk), .wr_en(wr_en), .addr(col), .data_in(r), .data_out(b0_out));
ram b1(.clk(clk), .wr_en(wr_en), .addr(col + 1), .data_in(b0_out), .data_out(b1_out));
ram b2(.clk(clk), .wr_en(wr_en), .addr(col + 2), .data_in(b1_out), .data_out(b2_out));
ram b3(.clk(clk), .wr_en(wr_en), .addr(col + 3), .data_in(b2_out), .data_out(b3_out));
ram b4(.clk(clk), .wr_en(wr_en), .addr(col + 4), .data_in(b3_out), .data_out(b4_out));
ram b5(.clk(clk), .wr_en(wr_en), .addr(col + 5), .data_in(b4_out), .data_out(b5_out));
ram b6(.clk(clk), .wr_en(wr_en), .addr(col + 6), .data_in(b5_out), .data_out(b6_out));
ram b7(.clk(clk), .wr_en(wr_en), .addr(col + 7), .data_in(b6_out), .data_out(b7_out));
ram b8(.clk(clk), .wr_en(wr_en), .addr(col + 8), .data_in(b7_out), .data_out(b8_out));
ram b9(.clk(clk), .wr_en(wr_en), .addr(col + 9), .data_in(b8_out), .data_out(b9_out));
ram b10(.clk(clk), .wr_en(wr_en), .addr(col + 10), .data_in(b9_out), .data_out(b10_out));

always @(*) begin




end
always @(posedge clk) begin

end

	initial begin 
	

	end

endmodule

module ram(
	input clk,
	input wr_en,
	input [9:0] addr, 
	input [7:0] data_in,
	output [7:0] data_out
);
	reg [7:0] mem [639:0] /* synthesis ramstyle = M10K */;
	initial begin
	mem[0] = 8'h00;
mem[1] = 8'h00;
mem[2] = 8'h00;
mem[3] = 8'h00;
mem[4] = 8'h00;
mem[5] = 8'h00;
mem[6] = 8'h00;
mem[7] = 8'h00;
mem[8] = 8'h00;
mem[9] = 8'h00;
mem[10] = 8'h00;
mem[11] = 8'h00;
mem[12] = 8'h00;
mem[13] = 8'h00;
mem[14] = 8'h00;
mem[15] = 8'h00;
mem[16] = 8'h00;
mem[17] = 8'h00;
mem[18] = 8'h00;
mem[19] = 8'h00;
mem[20] = 8'h00;
mem[21] = 8'h00;
mem[22] = 8'h00;
mem[23] = 8'h00;
mem[24] = 8'h00;
mem[25] = 8'h00;
mem[26] = 8'h00;
mem[27] = 8'h00;
mem[28] = 8'h00;
mem[29] = 8'h00;
mem[30] = 8'h00;
mem[31] = 8'h00;
mem[32] = 8'h00;
mem[33] = 8'h00;
mem[34] = 8'h00;
mem[35] = 8'h00;
mem[36] = 8'h00;
mem[37] = 8'h00;
mem[38] = 8'h00;
mem[39] = 8'h00;
mem[40] = 8'h00;
mem[41] = 8'h00;
mem[42] = 8'h00;
mem[43] = 8'h00;
mem[44] = 8'h00;
mem[45] = 8'h00;
mem[46] = 8'h00;
mem[47] = 8'h00;
mem[48] = 8'h00;
mem[49] = 8'h00;
mem[50] = 8'h00;
mem[51] = 8'h00;
mem[52] = 8'h00;
mem[53] = 8'h00;
mem[54] = 8'h00;
mem[55] = 8'h00;
mem[56] = 8'h00;
mem[57] = 8'h00;
mem[58] = 8'h00;
mem[59] = 8'h00;
mem[60] = 8'h00;
mem[61] = 8'h00;
mem[62] = 8'h00;
mem[63] = 8'h00;
mem[64] = 8'h00;
mem[65] = 8'h00;
mem[66] = 8'h00;
mem[67] = 8'h00;
mem[68] = 8'h00;
mem[69] = 8'h00;
mem[70] = 8'h00;
mem[71] = 8'h00;
mem[72] = 8'h00;
mem[73] = 8'h00;
mem[74] = 8'h00;
mem[75] = 8'h00;
mem[76] = 8'h00;
mem[77] = 8'h00;
mem[78] = 8'h00;
mem[79] = 8'h00;
mem[80] = 8'h00;
mem[81] = 8'h00;
mem[82] = 8'h00;
mem[83] = 8'h00;
mem[84] = 8'h00;
mem[85] = 8'h00;
mem[86] = 8'h00;
mem[87] = 8'h00;
mem[88] = 8'h00;
mem[89] = 8'h00;
mem[90] = 8'h00;
mem[91] = 8'h00;
mem[92] = 8'h00;
mem[93] = 8'h00;
mem[94] = 8'h00;
mem[95] = 8'h00;
mem[96] = 8'h00;
mem[97] = 8'h00;
mem[98] = 8'h00;
mem[99] = 8'h00;
mem[100] = 8'h00;
mem[101] = 8'h00;
mem[102] = 8'h00;
mem[103] = 8'h00;
mem[104] = 8'h00;
mem[105] = 8'h00;
mem[106] = 8'h00;
mem[107] = 8'h00;
mem[108] = 8'h00;
mem[109] = 8'h00;
mem[110] = 8'h00;
mem[111] = 8'h00;
mem[112] = 8'h00;
mem[113] = 8'h00;
mem[114] = 8'h00;
mem[115] = 8'h00;
mem[116] = 8'h00;
mem[117] = 8'h00;
mem[118] = 8'h00;
mem[119] = 8'h00;
mem[120] = 8'h00;
mem[121] = 8'h00;
mem[122] = 8'h00;
mem[123] = 8'h00;
mem[124] = 8'h00;
mem[125] = 8'h00;
mem[126] = 8'h00;
mem[127] = 8'h00;
mem[128] = 8'h00;
mem[129] = 8'h00;
mem[130] = 8'h00;
mem[131] = 8'h00;
mem[132] = 8'h00;
mem[133] = 8'h00;
mem[134] = 8'h00;
mem[135] = 8'h00;
mem[136] = 8'h00;
mem[137] = 8'h00;
mem[138] = 8'h00;
mem[139] = 8'h00;
mem[140] = 8'h00;
mem[141] = 8'h00;
mem[142] = 8'h00;
mem[143] = 8'h00;
mem[144] = 8'h00;
mem[145] = 8'h00;
mem[146] = 8'h00;
mem[147] = 8'h00;
mem[148] = 8'h00;
mem[149] = 8'h00;
mem[150] = 8'h00;
mem[151] = 8'h00;
mem[152] = 8'h00;
mem[153] = 8'h00;
mem[154] = 8'h00;
mem[155] = 8'h00;
mem[156] = 8'h00;
mem[157] = 8'h00;
mem[158] = 8'h00;
mem[159] = 8'h00;
mem[160] = 8'h00;
mem[161] = 8'h00;
mem[162] = 8'h00;
mem[163] = 8'h00;
mem[164] = 8'h00;
mem[165] = 8'h00;
mem[166] = 8'h00;
mem[167] = 8'h00;
mem[168] = 8'h00;
mem[169] = 8'h00;
mem[170] = 8'h00;
mem[171] = 8'h00;
mem[172] = 8'h00;
mem[173] = 8'h00;
mem[174] = 8'h00;
mem[175] = 8'h00;
mem[176] = 8'h00;
mem[177] = 8'h00;
mem[178] = 8'h00;
mem[179] = 8'h00;
mem[180] = 8'h00;
mem[181] = 8'h00;
mem[182] = 8'h00;
mem[183] = 8'h00;
mem[184] = 8'h00;
mem[185] = 8'h00;
mem[186] = 8'h00;
mem[187] = 8'h00;
mem[188] = 8'h00;
mem[189] = 8'h00;
mem[190] = 8'h00;
mem[191] = 8'h00;
mem[192] = 8'h00;
mem[193] = 8'h00;
mem[194] = 8'h00;
mem[195] = 8'h00;
mem[196] = 8'h00;
mem[197] = 8'h00;
mem[198] = 8'h00;
mem[199] = 8'h00;
mem[200] = 8'h00;
mem[201] = 8'h00;
mem[202] = 8'h00;
mem[203] = 8'h00;
mem[204] = 8'h00;
mem[205] = 8'h00;
mem[206] = 8'h00;
mem[207] = 8'h00;
mem[208] = 8'h00;
mem[209] = 8'h00;
mem[210] = 8'h00;
mem[211] = 8'h00;
mem[212] = 8'h00;
mem[213] = 8'h00;
mem[214] = 8'h00;
mem[215] = 8'h00;
mem[216] = 8'h00;
mem[217] = 8'h00;
mem[218] = 8'h00;
mem[219] = 8'h00;
mem[220] = 8'h00;
mem[221] = 8'h00;
mem[222] = 8'h00;
mem[223] = 8'h00;
mem[224] = 8'h00;
mem[225] = 8'h00;
mem[226] = 8'h00;
mem[227] = 8'h00;
mem[228] = 8'h00;
mem[229] = 8'h00;
mem[230] = 8'h00;
mem[231] = 8'h00;
mem[232] = 8'h00;
mem[233] = 8'h00;
mem[234] = 8'h00;
mem[235] = 8'h00;
mem[236] = 8'h00;
mem[237] = 8'h00;
mem[238] = 8'h00;
mem[239] = 8'h00;
mem[240] = 8'h00;
mem[241] = 8'h00;
mem[242] = 8'h00;
mem[243] = 8'h00;
mem[244] = 8'h00;
mem[245] = 8'h00;
mem[246] = 8'h00;
mem[247] = 8'h00;
mem[248] = 8'h00;
mem[249] = 8'h00;
mem[250] = 8'h00;
mem[251] = 8'h00;
mem[252] = 8'h00;
mem[253] = 8'h00;
mem[254] = 8'h00;
mem[255] = 8'h00;
mem[256] = 8'h00;
mem[257] = 8'h00;
mem[258] = 8'h00;
mem[259] = 8'h00;
mem[260] = 8'h00;
mem[261] = 8'h00;
mem[262] = 8'h00;
mem[263] = 8'h00;
mem[264] = 8'h00;
mem[265] = 8'h00;
mem[266] = 8'h00;
mem[267] = 8'h00;
mem[268] = 8'h00;
mem[269] = 8'h00;
mem[270] = 8'h00;
mem[271] = 8'h00;
mem[272] = 8'h00;
mem[273] = 8'h00;
mem[274] = 8'h00;
mem[275] = 8'h00;
mem[276] = 8'h00;
mem[277] = 8'h00;
mem[278] = 8'h00;
mem[279] = 8'h00;
mem[280] = 8'h00;
mem[281] = 8'h00;
mem[282] = 8'h00;
mem[283] = 8'h00;
mem[284] = 8'h00;
mem[285] = 8'h00;
mem[286] = 8'h00;
mem[287] = 8'h00;
mem[288] = 8'h00;
mem[289] = 8'h00;
mem[290] = 8'h00;
mem[291] = 8'h00;
mem[292] = 8'h00;
mem[293] = 8'h00;
mem[294] = 8'h00;
mem[295] = 8'h00;
mem[296] = 8'h00;
mem[297] = 8'h00;
mem[298] = 8'h00;
mem[299] = 8'h00;
mem[300] = 8'h00;
mem[301] = 8'h00;
mem[302] = 8'h00;
mem[303] = 8'h00;
mem[304] = 8'h00;
mem[305] = 8'h00;
mem[306] = 8'h00;
mem[307] = 8'h00;
mem[308] = 8'h00;
mem[309] = 8'h00;
mem[310] = 8'h00;
mem[311] = 8'h00;
mem[312] = 8'h00;
mem[313] = 8'h00;
mem[314] = 8'h00;
mem[315] = 8'h00;
mem[316] = 8'h00;
mem[317] = 8'h00;
mem[318] = 8'h00;
mem[319] = 8'h00;
mem[320] = 8'h00;
mem[321] = 8'h00;
mem[322] = 8'h00;
mem[323] = 8'h00;
mem[324] = 8'h00;
mem[325] = 8'h00;
mem[326] = 8'h00;
mem[327] = 8'h00;
mem[328] = 8'h00;
mem[329] = 8'h00;
mem[330] = 8'h00;
mem[331] = 8'h00;
mem[332] = 8'h00;
mem[333] = 8'h00;
mem[334] = 8'h00;
mem[335] = 8'h00;
mem[336] = 8'h00;
mem[337] = 8'h00;
mem[338] = 8'h00;
mem[339] = 8'h00;
mem[340] = 8'h00;
mem[341] = 8'h00;
mem[342] = 8'h00;
mem[343] = 8'h00;
mem[344] = 8'h00;
mem[345] = 8'h00;
mem[346] = 8'h00;
mem[347] = 8'h00;
mem[348] = 8'h00;
mem[349] = 8'h00;
mem[350] = 8'h00;
mem[351] = 8'h00;
mem[352] = 8'h00;
mem[353] = 8'h00;
mem[354] = 8'h00;
mem[355] = 8'h00;
mem[356] = 8'h00;
mem[357] = 8'h00;
mem[358] = 8'h00;
mem[359] = 8'h00;
mem[360] = 8'h00;
mem[361] = 8'h00;
mem[362] = 8'h00;
mem[363] = 8'h00;
mem[364] = 8'h00;
mem[365] = 8'h00;
mem[366] = 8'h00;
mem[367] = 8'h00;
mem[368] = 8'h00;
mem[369] = 8'h00;
mem[370] = 8'h00;
mem[371] = 8'h00;
mem[372] = 8'h00;
mem[373] = 8'h00;
mem[374] = 8'h00;
mem[375] = 8'h00;
mem[376] = 8'h00;
mem[377] = 8'h00;
mem[378] = 8'h00;
mem[379] = 8'h00;
mem[380] = 8'h00;
mem[381] = 8'h00;
mem[382] = 8'h00;
mem[383] = 8'h00;
mem[384] = 8'h00;
mem[385] = 8'h00;
mem[386] = 8'h00;
mem[387] = 8'h00;
mem[388] = 8'h00;
mem[389] = 8'h00;
mem[390] = 8'h00;
mem[391] = 8'h00;
mem[392] = 8'h00;
mem[393] = 8'h00;
mem[394] = 8'h00;
mem[395] = 8'h00;
mem[396] = 8'h00;
mem[397] = 8'h00;
mem[398] = 8'h00;
mem[399] = 8'h00;
mem[400] = 8'h00;
mem[401] = 8'h00;
mem[402] = 8'h00;
mem[403] = 8'h00;
mem[404] = 8'h00;
mem[405] = 8'h00;
mem[406] = 8'h00;
mem[407] = 8'h00;
mem[408] = 8'h00;
mem[409] = 8'h00;
mem[410] = 8'h00;
mem[411] = 8'h00;
mem[412] = 8'h00;
mem[413] = 8'h00;
mem[414] = 8'h00;
mem[415] = 8'h00;
mem[416] = 8'h00;
mem[417] = 8'h00;
mem[418] = 8'h00;
mem[419] = 8'h00;
mem[420] = 8'h00;
mem[421] = 8'h00;
mem[422] = 8'h00;
mem[423] = 8'h00;
mem[424] = 8'h00;
mem[425] = 8'h00;
mem[426] = 8'h00;
mem[427] = 8'h00;
mem[428] = 8'h00;
mem[429] = 8'h00;
mem[430] = 8'h00;
mem[431] = 8'h00;
mem[432] = 8'h00;
mem[433] = 8'h00;
mem[434] = 8'h00;
mem[435] = 8'h00;
mem[436] = 8'h00;
mem[437] = 8'h00;
mem[438] = 8'h00;
mem[439] = 8'h00;
mem[440] = 8'h00;
mem[441] = 8'h00;
mem[442] = 8'h00;
mem[443] = 8'h00;
mem[444] = 8'h00;
mem[445] = 8'h00;
mem[446] = 8'h00;
mem[447] = 8'h00;
mem[448] = 8'h00;
mem[449] = 8'h00;
mem[450] = 8'h00;
mem[451] = 8'h00;
mem[452] = 8'h00;
mem[453] = 8'h00;
mem[454] = 8'h00;
mem[455] = 8'h00;
mem[456] = 8'h00;
mem[457] = 8'h00;
mem[458] = 8'h00;
mem[459] = 8'h00;
mem[460] = 8'h00;
mem[461] = 8'h00;
mem[462] = 8'h00;
mem[463] = 8'h00;
mem[464] = 8'h00;
mem[465] = 8'h00;
mem[466] = 8'h00;
mem[467] = 8'h00;
mem[468] = 8'h00;
mem[469] = 8'h00;
mem[470] = 8'h00;
mem[471] = 8'h00;
mem[472] = 8'h00;
mem[473] = 8'h00;
mem[474] = 8'h00;
mem[475] = 8'h00;
mem[476] = 8'h00;
mem[477] = 8'h00;
mem[478] = 8'h00;
mem[479] = 8'h00;
mem[480] = 8'h00;
mem[481] = 8'h00;
mem[482] = 8'h00;
mem[483] = 8'h00;
mem[484] = 8'h00;
mem[485] = 8'h00;
mem[486] = 8'h00;
mem[487] = 8'h00;
mem[488] = 8'h00;
mem[489] = 8'h00;
mem[490] = 8'h00;
mem[491] = 8'h00;
mem[492] = 8'h00;
mem[493] = 8'h00;
mem[494] = 8'h00;
mem[495] = 8'h00;
mem[496] = 8'h00;
mem[497] = 8'h00;
mem[498] = 8'h00;
mem[499] = 8'h00;
mem[500] = 8'h00;
mem[501] = 8'h00;
mem[502] = 8'h00;
mem[503] = 8'h00;
mem[504] = 8'h00;
mem[505] = 8'h00;
mem[506] = 8'h00;
mem[507] = 8'h00;
mem[508] = 8'h00;
mem[509] = 8'h00;
mem[510] = 8'h00;
mem[511] = 8'h00;
mem[512] = 8'h00;
mem[513] = 8'h00;
mem[514] = 8'h00;
mem[515] = 8'h00;
mem[516] = 8'h00;
mem[517] = 8'h00;
mem[518] = 8'h00;
mem[519] = 8'h00;
mem[520] = 8'h00;
mem[521] = 8'h00;
mem[522] = 8'h00;
mem[523] = 8'h00;
mem[524] = 8'h00;
mem[525] = 8'h00;
mem[526] = 8'h00;
mem[527] = 8'h00;
mem[528] = 8'h00;
mem[529] = 8'h00;
mem[530] = 8'h00;
mem[531] = 8'h00;
mem[532] = 8'h00;
mem[533] = 8'h00;
mem[534] = 8'h00;
mem[535] = 8'h00;
mem[536] = 8'h00;
mem[537] = 8'h00;
mem[538] = 8'h00;
mem[539] = 8'h00;
mem[540] = 8'h00;
mem[541] = 8'h00;
mem[542] = 8'h00;
mem[543] = 8'h00;
mem[544] = 8'h00;
mem[545] = 8'h00;
mem[546] = 8'h00;
mem[547] = 8'h00;
mem[548] = 8'h00;
mem[549] = 8'h00;
mem[550] = 8'h00;
mem[551] = 8'h00;
mem[552] = 8'h00;
mem[553] = 8'h00;
mem[554] = 8'h00;
mem[555] = 8'h00;
mem[556] = 8'h00;
mem[557] = 8'h00;
mem[558] = 8'h00;
mem[559] = 8'h00;
mem[560] = 8'h00;
mem[561] = 8'h00;
mem[562] = 8'h00;
mem[563] = 8'h00;
mem[564] = 8'h00;
mem[565] = 8'h00;
mem[566] = 8'h00;
mem[567] = 8'h00;
mem[568] = 8'h00;
mem[569] = 8'h00;
mem[570] = 8'h00;
mem[571] = 8'h00;
mem[572] = 8'h00;
mem[573] = 8'h00;
mem[574] = 8'h00;
mem[575] = 8'h00;
mem[576] = 8'h00;
mem[577] = 8'h00;
mem[578] = 8'h00;
mem[579] = 8'h00;
mem[580] = 8'h00;
mem[581] = 8'h00;
mem[582] = 8'h00;
mem[583] = 8'h00;
mem[584] = 8'h00;
mem[585] = 8'h00;
mem[586] = 8'h00;
mem[587] = 8'h00;
mem[588] = 8'h00;
mem[589] = 8'h00;
mem[590] = 8'h00;
mem[591] = 8'h00;
mem[592] = 8'h00;
mem[593] = 8'h00;
mem[594] = 8'h00;
mem[595] = 8'h00;
mem[596] = 8'h00;
mem[597] = 8'h00;
mem[598] = 8'h00;
mem[599] = 8'h00;
mem[600] = 8'h00;
mem[601] = 8'h00;
mem[602] = 8'h00;
mem[603] = 8'h00;
mem[604] = 8'h00;
mem[605] = 8'h00;
mem[606] = 8'h00;
mem[607] = 8'h00;
mem[608] = 8'h00;
mem[609] = 8'h00;
mem[610] = 8'h00;
mem[611] = 8'h00;
mem[612] = 8'h00;
mem[613] = 8'h00;
mem[614] = 8'h00;
mem[615] = 8'h00;
mem[616] = 8'h00;
mem[617] = 8'h00;
mem[618] = 8'h00;
mem[619] = 8'h00;
mem[620] = 8'h00;
mem[621] = 8'h00;
mem[622] = 8'h00;
mem[623] = 8'h00;
mem[624] = 8'h00;
mem[625] = 8'h00;
mem[626] = 8'h00;
mem[627] = 8'h00;
mem[628] = 8'h00;
mem[629] = 8'h00;
mem[630] = 8'h00;
mem[631] = 8'h00;
mem[632] = 8'h00;
mem[633] = 8'h00;
mem[634] = 8'h00;
mem[635] = 8'h00;
mem[636] = 8'h00;
mem[637] = 8'h00;
mem[638] = 8'h00;
mem[639] = 8'h00;
	end
	always @(posedge clk) begin
		if(wr_en == 1'b1) begin
			mem[addr] <= #1 data_in;
		end
	end
	assign data_out = mem[addr];
endmodule

