module gauss(
input clk,
input [7:0] r, b , g,
input [12:0] col,
input buff_en,
input shift_en,
input [1:0] filt_sel,
output reg [7:0] out_r, out_g, out_b

);

reg [1:0] k_sel;
reg [20:0] tmp_1[2:0]; 
reg [7:0] buff [639:0] [2:0];
reg [7:0] shift [10:0] [639:0] [2:0];
saturate satr(.in(tmp_1[0][17:8]), .out(out_r));
saturate satb(.in(tmp_1[1][17:8]), .out(out_g));
saturate satg(.in(tmp_1[2][17:8]), .out(out_b));
wire [7:0] gauss_r, gauss_g, gauss_b;

integer color, column;
integer temp1, temp2, temp3, temp4;
reg [7:0] mem[10:0][10:0][2:0];

always @(*) begin
	
	case(filt_sel)
		2'b01: begin
			k_sel = 2'b00;
		end
		2'b10: begin
			k_sel = 2'b01;
		end
		default begin
			k_sel = 2'b10;
		end
	
	endcase
end
always @(posedge clk) begin
	for(temp3 = 0; temp3 <= 2; temp3 = temp3 + 1) begin
		tmp_1[temp3] = 21'b0;
		for(temp2 = 0; temp2 <= 4; temp2 = temp2 + 1) begin
			tmp_1[temp3] = tmp_1[temp3] + 
						mem[temp2][10][k_sel] * shift[10][col + 5][temp3] + 
						mem[temp2][9][k_sel] * shift[10][col + 4][temp3] + 
						mem[temp2][8][k_sel] * shift[10][col + 3][temp3] + 
						mem[temp2][7][k_sel] * shift[10][col + 2][temp3] + 
						mem[temp2][6][k_sel] * shift[10][col + 1][temp3] +
						mem[temp2][5][k_sel] * shift[10][col][temp3] 	 + 
						mem[temp2][4][k_sel] * shift[10][col - 1][temp3] + 
						mem[temp2][3][k_sel] * shift[10][col - 2][temp3] + 
						mem[temp2][2][k_sel] * shift[10][col - 3][temp3] + 
						mem[temp2][1][k_sel] * shift[10][col - 4][temp3] +
						mem[temp2][0][k_sel] * shift[10][col - 5][temp3];
		end
	end

//	for(temp4 = 0; temp4 <= 2; temp4 = temp4 + 1)begin
//		tmp_2[temp4] = (tmp_1[temp4] * 8'b0000101);
//	end

//	8'b00000100 * shift[9][col - 2][0] + 
//	8'b00001111 * shift[9][col - 1][0] + 
//	8'b00011000 * shift[9][col][0] + 
//	8'b00001111 * shift[9][col + 1][0] + 
//	8'b00000100 * shift[9][col + 2][0] + 
//	8'b00000110 * shift[8][col - 2][0] + 
//	8'b00011000 * shift[8][col - 1][0] + 
//	8'b00100110 * shift[8][col][0] + 
//	8'b00011000 * shift[8][col + 1][0] + 
//	8'b00000110 * shift[8][col + 2][0] + 
//	8'b00000100 * shift[7][col - 2][0] + 
//	8'b00001111 * shift[7][col - 1][0] + 
//	8'b00011000 * shift[7][col][0] + 
//	8'b00001111 * shift[7][col + 1][0] + 
//	8'b00000100 * shift[7][col + 2][0] + 
//	8'b00000001 * shift[6][col - 2][0] + 
//	8'b00000100 * shift[6][col - 1][0] + 
//	8'b00000110 * shift[6][col][0] + 
//	8'b00000100 * shift[6][col + 1][0] + 
//	8'b00000001 * shift[6][col + 2][0];
//	tmp_g1 = 8'b00000001 * shift[10][col - 2][1] + 
//	8'b00000100 * shift[10][col - 1][1] + 
//	8'b00000110 * shift[10][col][1] + 
//	8'b00000100 * shift[10][col + 1][1] + 
//	8'b00000001 * shift[10][col + 2][1] + 
//	8'b00000100 * shift[9][col - 2][1] + 
//	8'b00001111 * shift[9][col - 1][1] + 
//	8'b00011000 * shift[9][col][1] + 
//	8'b00001111 * shift[9][col + 1][1] + 
//	8'b00000100 * shift[9][col + 2][1] + 
//	8'b00000110 * shift[8][col - 2][1] + 
//	8'b00011000 * shift[8][col - 1][1] + 
//	8'b00100110 * shift[8][col][1] + 
//	8'b00011000 * shift[8][col + 1][1] + 
//	8'b00000110 * shift[8][col + 2][1] + 
//	8'b00000100 * shift[7][col - 2][1] + 
//	8'b00001111 * shift[7][col - 1][1] + 
//	8'b00011000 * shift[7][col][1] + 
//	8'b00001111 * shift[7][col + 1][1] + 
//	8'b00000100 * shift[7][col + 2][1] + 
//	8'b00000001 * shift[6][col - 2][1] + 
//	8'b00000100 * shift[6][col - 1][1] + 
//	8'b00000110 * shift[6][col][1] + 
//	8'b00000100 * shift[6][col + 1][1] + 
//	8'b00000001 * shift[6][col + 2][1];
//	tmp_g2 = (tmp_g1 * 8'b0000101);
//	tmp_b1 = 8'b00000001 * shift[10][col - 2][2] + 
//	8'b00000100 * shift[10][col - 1][2] + 
//	8'b00000110 * shift[10][col][2] + 
//	8'b00000100 * shift[10][col + 1][2] + 
//	8'b00000001 * shift[10][col + 2][2] + 
//	8'b00000100 * shift[9][col - 2][2] + 
//	8'b00001111 * shift[9][col - 1][2] + 
//	8'b00011000 * shift[9][col][2] + 
//	8'b00001111 * shift[9][col + 1][2] + 
//	8'b00000100 * shift[9][col + 2][2] + 
//	8'b00000110 * shift[8][col - 2][2] + 
//	8'b00011000 * shift[8][col - 1][2] + 
//	8'b00100110 * shift[8][col][2] + 
//	8'b00011000 * shift[8][col + 1][2] + 
//	8'b00000110 * shift[8][col + 2][2] + 
//	8'b00000100 * shift[7][col - 2][2] + 
//	8'b00001111 * shift[7][col - 1][2] + 
//	8'b00011000 * shift[7][col][2] + 
//	8'b00001111 * shift[7][col + 1][2] + 
//	8'b00000100 * shift[7][col + 2][2] + 
//	8'b00000001 * shift[6][col - 2][2] + 
//	8'b00000100 * shift[6][col - 1][2] + 
//	8'b00000110 * shift[6][col][2] + 
//	8'b00000100 * shift[6][col + 1][2] + 
//	8'b00000001 * shift[6][col + 2][2];
//	tmp_b2 = (tmp_b1 * 8'b0000101);

end
always @(posedge clk) begin
	if( buff_en == 1'b1) begin
		buff[col][0] <= #1 r;
		buff[col][1] <= #1 g;
		buff[col][2] <= #1 b;
	end
	if(shift_en == 1'b1) begin
		for(color = 0; color < 3; color = color + 1)begin
			for(column = 0; column < 640; column = column + 1) begin
				shift[0][column][color] <= #1 buff[column][color];
				shift[1][column][color] <= #1 shift[0][column][color];
				shift[2][column][color] <= #1 shift[1][column][color];
				shift[3][column][color] <= #1 shift[2][column][color];
				shift[4][column][color] <= #1 shift[3][column][color];
				shift[5][column][color] <= #1 shift[4][column][color];
				shift[6][column][color] <= #1 shift[5][column][color];
				shift[7][column][color] <= #1 shift[6][column][color];
				shift[8][column][color] <= #1 shift[7][column][color];
				shift[9][column][color] <= #1 shift[8][column][color];
				shift[10][column][color] <= #1 shift[9][column][color];
			end
		end
	end
	
end

	initial begin 
		mem[0][0][0] = 8'b00000000;
		mem[0][0][1] = 8'b00000001;
		mem[0][1][0] = 8'b00000000;
		mem[0][1][1] = 8'b00000001;
		mem[0][2][0] = 8'b00000000;
		mem[0][2][1] = 8'b00000010;
		mem[0][3][0] = 8'b00000000;
		mem[0][3][1] = 8'b00000010;
		mem[0][4][0] = 8'b00000000;
		mem[0][4][1] = 8'b00000010;
		mem[0][5][0] = 8'b00000000;
		mem[0][5][1] = 8'b00000010;
		mem[0][6][0] = 8'b00000000;
		mem[0][6][1] = 8'b00000010;
		mem[0][7][0] = 8'b00000000;
		mem[0][7][1] = 8'b00000010;
		mem[0][8][0] = 8'b00000000;
		mem[0][8][1] = 8'b00000010;
		mem[0][9][0] = 8'b00000000;
		mem[0][9][1] = 8'b00000001;
		mem[0][10][0] = 8'b00000000;
		mem[0][10][1] = 8'b00000001;
		mem[1][0][0] = 8'b00000000;
		mem[1][0][1] = 8'b00000001;
		mem[1][1][0] = 8'b00000000;
		mem[1][1][1] = 8'b00000010;
		mem[1][2][0] = 8'b00000000;
		mem[1][2][1] = 8'b00000010;
		mem[1][3][0] = 8'b00000000;
		mem[1][3][1] = 8'b00000010;
		mem[1][4][0] = 8'b00000000;
		mem[1][4][1] = 8'b00000010;
		mem[1][5][0] = 8'b00000000;
		mem[1][5][1] = 8'b00000010;
		mem[1][6][0] = 8'b00000000;
		mem[1][6][1] = 8'b00000010;
		mem[1][7][0] = 8'b00000000;
		mem[1][7][1] = 8'b00000010;
		mem[1][8][0] = 8'b00000000;
		mem[1][8][1] = 8'b00000010;
		mem[1][9][0] = 8'b00000000;
		mem[1][9][1] = 8'b00000010;
		mem[1][10][0] = 8'b00000000;
		mem[1][10][1] = 8'b00000001;
		mem[2][0][0] = 8'b00000000;
		mem[2][0][1] = 8'b00000010;
		mem[2][1][0] = 8'b00000000;
		mem[2][1][1] = 8'b00000010;
		mem[2][2][0] = 8'b00000000;
		mem[2][2][1] = 8'b00000010;
		mem[2][3][0] = 8'b00000000;
		mem[2][3][1] = 8'b00000010;
		mem[2][4][0] = 8'b00000000;
		mem[2][4][1] = 8'b00000011;
		mem[2][5][0] = 8'b00000000;
		mem[2][5][1] = 8'b00000011;
		mem[2][6][0] = 8'b00000000;
		mem[2][6][1] = 8'b00000011;
		mem[2][7][0] = 8'b00000000;
		mem[2][7][1] = 8'b00000010;
		mem[2][8][0] = 8'b00000000;
		mem[2][8][1] = 8'b00000010;
		mem[2][9][0] = 8'b00000000;
		mem[2][9][1] = 8'b00000010;
		mem[2][10][0] = 8'b00000000;
		mem[2][10][1] = 8'b00000010;
		mem[3][0][0] = 8'b00000000;
		mem[3][0][1] = 8'b00000010;
		mem[3][1][0] = 8'b00000000;
		mem[3][1][1] = 8'b00000010;
		mem[3][2][0] = 8'b00000000;
		mem[3][2][1] = 8'b00000010;
		mem[3][3][0] = 8'b00001001;
		mem[3][3][1] = 8'b00000011;
		mem[3][4][0] = 8'b00001010;
		mem[3][4][1] = 8'b00000011;
		mem[3][5][0] = 8'b00001010;
		mem[3][5][1] = 8'b00000011;
		mem[3][6][0] = 8'b00001010;
		mem[3][6][1] = 8'b00000011;
		mem[3][7][0] = 8'b00001001;
		mem[3][7][1] = 8'b00000011;
		mem[3][8][0] = 8'b00000000;
		mem[3][8][1] = 8'b00000010;
		mem[3][9][0] = 8'b00000000;
		mem[3][9][1] = 8'b00000010;
		mem[3][10][0] = 8'b00000000;
		mem[3][10][1] = 8'b00000010;
		mem[4][0][0] = 8'b00000000;
		mem[4][0][1] = 8'b00000010;
		mem[4][1][0] = 8'b00000000;
		mem[4][1][1] = 8'b00000010;
		mem[4][2][0] = 8'b00000000;
		mem[4][2][1] = 8'b00000011;
		mem[4][3][0] = 8'b00001010;
		mem[4][3][1] = 8'b00000011;
		mem[4][4][0] = 8'b00001011;
		mem[4][4][1] = 8'b00000011;
		mem[4][5][0] = 8'b00001011;
		mem[4][5][1] = 8'b00000011;
		mem[4][6][0] = 8'b00001011;
		mem[4][6][1] = 8'b00000011;
		mem[4][7][0] = 8'b00001010;
		mem[4][7][1] = 8'b00000011;
		mem[4][8][0] = 8'b00000000;
		mem[4][8][1] = 8'b00000011;
		mem[4][9][0] = 8'b00000000;
		mem[4][9][1] = 8'b00000010;
		mem[4][10][0] = 8'b00000000;
		mem[4][10][1] = 8'b00000010;
		mem[5][0][0] = 8'b00000000;
		mem[5][0][1] = 8'b00000010;
		mem[5][1][0] = 8'b00000000;
		mem[5][1][1] = 8'b00000010;
		mem[5][2][0] = 8'b00000000;
		mem[5][2][1] = 8'b00000011;
		mem[5][3][0] = 8'b00001010;
		mem[5][3][1] = 8'b00000011;
		mem[5][4][0] = 8'b00001011;
		mem[5][4][1] = 8'b00000011;
		mem[5][5][0] = 8'b00001011;
		mem[5][5][1] = 8'b00000011;
		mem[5][6][0] = 8'b00001011;
		mem[5][6][1] = 8'b00000011;
		mem[5][7][0] = 8'b00001010;
		mem[5][7][1] = 8'b00000011;
		mem[5][8][0] = 8'b00000000;
		mem[5][8][1] = 8'b00000011;
		mem[5][9][0] = 8'b00000000;
		mem[5][9][1] = 8'b00000010;
		mem[5][10][0] = 8'b00000000;
		mem[5][10][1] = 8'b00000010;
		mem[6][0][0] = 8'b00000000;
		mem[6][0][1] = 8'b00000010;
		mem[6][1][0] = 8'b00000000;
		mem[6][1][1] = 8'b00000010;
		mem[6][2][0] = 8'b00000000;
		mem[6][2][1] = 8'b00000011;
		mem[6][3][0] = 8'b00001010;
		mem[6][3][1] = 8'b00000011;
		mem[6][4][0] = 8'b00001011;
		mem[6][4][1] = 8'b00000011;
		mem[6][5][0] = 8'b00001011;
		mem[6][5][1] = 8'b00000011;
		mem[6][6][0] = 8'b00001011;
		mem[6][6][1] = 8'b00000011;
		mem[6][7][0] = 8'b00001010;
		mem[6][7][1] = 8'b00000011;
		mem[6][8][0] = 8'b00000000;
		mem[6][8][1] = 8'b00000011;
		mem[6][9][0] = 8'b00000000;
		mem[6][9][1] = 8'b00000010;
		mem[6][10][0] = 8'b00000000;
		mem[6][10][1] = 8'b00000010;
		mem[7][0][0] = 8'b00000000;
		mem[7][0][1] = 8'b00000010;
		mem[7][1][0] = 8'b00000000;
		mem[7][1][1] = 8'b00000010;
		mem[7][2][0] = 8'b00000000;
		mem[7][2][1] = 8'b00000010;
		mem[7][3][0] = 8'b00001001;
		mem[7][3][1] = 8'b00000011;
		mem[7][4][0] = 8'b00001010;
		mem[7][4][1] = 8'b00000011;
		mem[7][5][0] = 8'b00001010;
		mem[7][5][1] = 8'b00000011;
		mem[7][6][0] = 8'b00001010;
		mem[7][6][1] = 8'b00000011;
		mem[7][7][0] = 8'b00001001;
		mem[7][7][1] = 8'b00000011;
		mem[7][8][0] = 8'b00000000;
		mem[7][8][1] = 8'b00000010;
		mem[7][9][0] = 8'b00000000;
		mem[7][9][1] = 8'b00000010;
		mem[7][10][0] = 8'b00000000;
		mem[7][10][1] = 8'b00000010;
		mem[8][0][0] = 8'b00000000;
		mem[8][0][1] = 8'b00000010;
		mem[8][1][0] = 8'b00000000;
		mem[8][1][1] = 8'b00000010;
		mem[8][2][0] = 8'b00000000;
		mem[8][2][1] = 8'b00000010;
		mem[8][3][0] = 8'b00000000;
		mem[8][3][1] = 8'b00000010;
		mem[8][4][0] = 8'b00000000;
		mem[8][4][1] = 8'b00000011;
		mem[8][5][0] = 8'b00000000;
		mem[8][5][1] = 8'b00000011;
		mem[8][6][0] = 8'b00000000;
		mem[8][6][1] = 8'b00000011;
		mem[8][7][0] = 8'b00000000;
		mem[8][7][1] = 8'b00000010;
		mem[8][8][0] = 8'b00000000;
		mem[8][8][1] = 8'b00000010;
		mem[8][9][0] = 8'b00000000;
		mem[8][9][1] = 8'b00000010;
		mem[8][10][0] = 8'b00000000;
		mem[8][10][1] = 8'b00000010;
		mem[9][0][0] = 8'b00000000;
		mem[9][0][1] = 8'b00000001;
		mem[9][1][0] = 8'b00000000;
		mem[9][1][1] = 8'b00000010;
		mem[9][2][0] = 8'b00000000;
		mem[9][2][1] = 8'b00000010;
		mem[9][3][0] = 8'b00000000;
		mem[9][3][1] = 8'b00000010;
		mem[9][4][0] = 8'b00000000;
		mem[9][4][1] = 8'b00000010;
		mem[9][5][0] = 8'b00000000;
		mem[9][5][1] = 8'b00000010;
		mem[9][6][0] = 8'b00000000;
		mem[9][6][1] = 8'b00000010;
		mem[9][7][0] = 8'b00000000;
		mem[9][7][1] = 8'b00000010;
		mem[9][8][0] = 8'b00000000;
		mem[9][8][1] = 8'b00000010;
		mem[9][9][0] = 8'b00000000;
		mem[9][9][1] = 8'b00000010;
		mem[9][10][0] = 8'b00000000;
		mem[9][10][1] = 8'b00000001;
		mem[10][0][0] = 8'b00000000;
		mem[10][0][1] = 8'b00000001;
		mem[10][1][0] = 8'b00000000;
		mem[10][1][1] = 8'b00000001;
		mem[10][2][0] = 8'b00000000;
		mem[10][2][1] = 8'b00000010;
		mem[10][3][0] = 8'b00000000;
		mem[10][3][1] = 8'b00000010;
		mem[10][4][0] = 8'b00000000;
		mem[10][4][1] = 8'b00000010;
		mem[10][5][0] = 8'b00000000;
		mem[10][5][1] = 8'b00000010;
		mem[10][6][0] = 8'b00000000;
		mem[10][6][1] = 8'b00000010;
		mem[10][7][0] = 8'b00000000;
		mem[10][7][1] = 8'b00000010;
		mem[10][8][0] = 8'b00000000;
		mem[10][8][1] = 8'b00000010;
		mem[10][9][0] = 8'b00000000;
		mem[10][9][1] = 8'b00000001;
		mem[10][10][0] = 8'b00000000;
		mem[10][10][1] = 8'b00000001;
		integer mem2, mem3;
		for(mem2 = 0; mem < 11; mem2 = mem2 + 1) begin
			for(mem3 = 0; mem3 < 11; mem3 = mem3 + 1)begin
				if(mem2 == 3'd5 && mem3 == 3'd5)begin
					mem[mem2][mem3][2] = 8'b1111_1111;
				end
				else mem[mem2][mem3][2] = 8'b0000_0000;

			end
		end
	end
	

endmodule

